// simple_cpu.v - Top-level module for the Simple CPU on DE10-Standard

module simple_cpu (
    input wire clk_50mhz,    // 50MHz clock from DE10-Standard
    input wire key0_n,       // Active-low reset button (KEY0)
    // 偵錯輸出埠：方便 ModelSim 觀察內部訊號，或未來連接到 FPGA LED
    output wire [7:0] debug_output_acc,      // 顯示累加器內容
    output wire [7:0] debug_pc_out,          // 顯示 PC 值
    output wire [15:0] debug_instruction_out // 顯示當前指令
);

    // --- Define Instruction Opcodes for top-level use ---
    // These must match the parameter definitions in ir_decoder.v
    parameter OP_NO_OP          = 8'h00;
    parameter OP_LOAD_ACC_IMM   = 8'h10;
    parameter OP_LOAD_ACC_MEM   = 8'h11;
    parameter OP_STORE_ACC_MEM  = 8'h20;
    parameter OP_ADD_ACC_IMM    = 8'h30;
    parameter OP_ADD_ACC_MEM    = 8'h31;
    parameter OP_SUB_ACC_IMM    = 8'h40;
    parameter OP_SUB_ACC_MEM    = 8'h41;
    parameter OP_AND_ACC_IMM    = 8'h50;
    parameter OP_AND_ACC_MEM    = 8'h51;
    parameter OP_INC_ACC        = 8'h60;
    parameter OP_JUMP           = 8'h70;
    parameter OP_OUT_ACC_SERIAL = 8'h80;


    // --- Internal Wires and Registers ---

    // PC related signals
    wire [7:0] pc_out;
    wire pc_load_en;
    wire [7:0] jump_addr;

    // RAM related signals
    wire [7:0] ram_addr;                 // Address for RAM access (PC or Operand)
    wire [15:0] instruction_from_ram;    // 16-bit instruction/data fetched from RAM
    wire ram_we;                         // RAM Write Enable
    wire [15:0] ram_data_in;             // Data to write to RAM (from ACC for STORE)

    // IR Decoder related signals (control signals generated by decoder)
    wire [7:0] decoded_immediate_operand; // 8-bit operand from instruction
    wire ram_addr_mux_sel;               // Mux select for RAM address (0: PC, 1: Operand)
    wire [3:0] alu_opcode;
    wire alu_a_mux_sel;                  // Not strictly used, ALU A is always ACC
    wire alu_b_mux_sel;                  // Select for ALU B (Immediate or RAM_data_out_lower8bits)
    wire acc_load_en;                    // Accumulator load enable
    wire serial_out_en;                  // 內部訊號：來自 ir_decoder，但不再連接到外部 UART 硬體
    wire [7:0] decoded_opcode;           // Wire to connect to ir_decoder's decoded_opcode_out

    // ACC related signals
    wire [7:0] acc_out;
    wire [7:0] acc_data_in_muxed;        // Data routed to ACC for loading

    // ALU related signals
    wire [7:0] alu_a_input;
    wire [7:0] alu_b_input;
    wire [7:0] alu_result;
    wire alu_carry_out;                  // ALU carry out flag

    // --- Component Instantiations ---

    // 1. Program Counter
    program_counter u_pc (
        .clk(clk_50mhz),
        .reset_n(key0_n),
        .load_en(pc_load_en),
        .next_addr_in(jump_addr),
        .pc_out(pc_out)
    );

    // 2. RAM (Instruction & Data Memory) - 使用 IP Catalog 生成的模組
    // 根據 ram_inst.txt (ram_inst.v) 提供的埠名稱與 simple_cpu 訊號對應
    ram u_ram ( // 模組名稱是 ram，實例名稱為 u_ram
        .address ( ram_addr ),               // IP Port: .address  <-- 連接 simple_cpu 的 ram_addr
        .clock   ( clk_50mhz ),              // IP Port: .clock    <-- 連接 simple_cpu 的 clk_50mhz
        .data    ( ram_data_in ),            // IP Port: .data     <-- 連接 simple_cpu 的 ram_data_in
        .wren    ( ram_we ),                 // IP Port: .wren     <-- 連接 simple_cpu 的 ram_we
        .q       ( instruction_from_ram )    // IP Port: .q        <-- 連接 simple_cpu 的 instruction_from_ram
    );

    // Mux for RAM Address: Selects between PC (for instruction fetch) and Operand (for data access)
    assign ram_addr = (ram_addr_mux_sel == 1'b1) ? decoded_immediate_operand : pc_out;

    // Data to write to RAM for STORE instruction: Comes from Accumulator
    assign ram_data_in = {8'h00, acc_out};

    // 3. Instruction Register (IR) / Decoder
    ir_decoder u_ir_decoder (
        .clk(clk_50mhz),
        .reset_n(key0_n),
        .instruction_in(instruction_from_ram),

        .pc_load_en(pc_load_en),
        .jump_addr(jump_addr),

        .ram_we(ram_we),
        .ram_addr_mux_sel(ram_addr_mux_sel),

        .alu_opcode(alu_opcode),
        .alu_a_mux_sel(alu_a_mux_sel),
        .alu_b_mux_sel(alu_b_mux_sel),

        .acc_load_en(acc_load_en),

        .immediate_operand(decoded_immediate_operand),
        .serial_out_en(serial_out_en), // serial_out_en 作為內部連接線
        .decoded_opcode_out(decoded_opcode)
    );

    // 4. Accumulator
    accumulator u_acc (
        .clk(clk_50mhz),
        .reset_n(key0_n),
        .acc_load_en(acc_load_en),
        .data_in(acc_data_in_muxed),
        .acc_out(acc_out)
    );

    // Mux for Accumulator Data Input: Selects source for ACC loading
    assign acc_data_in_muxed =
        (decoded_opcode == OP_LOAD_ACC_IMM)  ? decoded_immediate_operand :
        (decoded_opcode == OP_LOAD_ACC_MEM)  ? instruction_from_ram[7:0] :
        alu_result;

    // 5. ALU
    alu u_alu (
        .a(alu_a_input),
        .b(alu_b_input),
        .opcode(alu_opcode),
        .result(alu_result),
        .carry_out(alu_carry_out)
    );

    // Mux for ALU Operand A: In this simple CPU, ALU A is always from Accumulator
    assign alu_a_input = acc_out;

    // Mux for ALU Operand B: Selects between Immediate_Operand and Lower 8 bits of RAM data
    assign alu_b_input = (alu_b_mux_sel == 1'b0) ? decoded_immediate_operand : instruction_from_ram[7:0];

    // --- 偵錯輸出連接 ---
    assign debug_output_acc = acc_out;
    assign debug_pc_out = pc_out;
    assign debug_instruction_out = instruction_from_ram;

endmodule