// simple_cpu.v - Top-level module for the Simple CPU on DE10-Standard

module simple_cpu (
    input wire clk_50mhz,        // 50MHz clock from DE10-Standard
    input wire key0_n,            // Active-low reset button (KEY0)
    // 偵錯輸出埠：方便 ModelSim 觀察內部訊號，或未來連接到 FPGA LED
    output wire [7:0] debug_output_acc,      // 顯示累加器內容
    output wire [7:0] debug_pc_out,          // 顯示 PC 值
    output wire [15:0] debug_instruction_out // 顯示當前指令
);

    // --- Define Instruction Opcodes for top-level use ---
    // These must match the parameter definitions in ir_decoder.v
    parameter OP_NO_OP            = 8'h00;
    parameter OP_LOAD_ACC_IMM     = 8'h10;
    parameter OP_LOAD_ACC_MEM     = 8'h11;
    parameter OP_STORE_ACC_MEM    = 8'h20;
    parameter OP_ADD_ACC_IMM      = 8'h30;
    parameter OP_ADD_ACC_MEM      = 8'h31;
    parameter OP_SUB_ACC_IMM      = 8'h40;
    parameter OP_SUB_ACC_MEM      = 8'h41;
    parameter OP_AND_ACC_IMM      = 8'h50;
    parameter OP_AND_ACC_MEM      = 8'h51;
    parameter OP_INC_ACC          = 8'h60;
    parameter OP_JUMP             = 8'h70;
    parameter OP_OUT_ACC_SERIAL   = 8'h80;


    // --- Internal Wires and Registers ---

    // PC related signals
    wire [7:0] pc_out;
    wire pc_load_en;
    wire [7:0] jump_addr;

    // RAM related signals (Now using two ports)
    // Port A: Instruction Fetch
    wire [15:0] instruction_from_ram_inst; // 16-bit instruction fetched from RAM (Port A)

    // Port B: Data Access
    wire [7:0] ram_data_addr;           // Address for RAM data access (Operand)
    wire [15:0] ram_data_in_data;       // Data to write to RAM (from ACC for STORE)
    wire ram_we_data;                   // RAM Write Enable for data port
    wire [15:0] data_from_ram_data;     // 16-bit data fetched from RAM (Port B)


    // IR Decoder related signals (control signals generated by decoder)
    wire [7:0] decoded_immediate_operand; // 8-bit operand from instruction
    // wire ram_addr_mux_sel;             // NO LONGER NEEDED with dual-port RAM for address muxing
    wire [3:0] alu_opcode;
    wire alu_a_mux_sel;                  // Not strictly used, ALU A is always ACC
    wire alu_b_mux_sel;                  // Select for ALU B (Immediate or RAM_data_out_lower8bits)
    wire acc_load_en;                    // Accumulator load enable
    wire serial_out_en;                  // 內部訊號：來自 ir_decoder
    wire [7:0] decoded_opcode;           // Wire to connect to ir_decoder's decoded_opcode_out

    // ACC related signals
    wire [7:0] acc_out;
    wire [7:0] acc_data_in_muxed;        // Data routed to ACC for loading

    // ALU related signals
    wire [7:0] alu_a_input;
    wire [7:0] alu_b_input;
    wire [7:0] alu_result;
    wire alu_carry_out;                  // ALU carry out flag

    // --- Component Instantiations ---

    // 1. Program Counter
    program_counter u_pc (
        .clk(clk_50mhz),
        .reset_n(key0_n),
        .load_en(pc_load_en),
        .next_addr_in(jump_addr),
        .pc_out(pc_out)
    );

    // 2. RAM (Instruction & Data Memory) - NOW DUAL-PORT RAM
    ram u_ram (
        .clk(clk_50mhz),

        // Port A: Instruction Fetch
        .addr_a(pc_out),                        // PC directly feeds instruction address
        .data_out_a(instruction_from_ram_inst), // Instruction comes out from this port

        // Port B: Data Access
        .we_b(ram_we_data),                     // Write Enable from IR Decoder
        .addr_b(ram_data_addr),                 // Data address from IR Decoder (Operand)
        .data_in_b(ram_data_in_data),           // Data to write (from ACC)
        .data_out_b(data_from_ram_data)         // Data read from memory
    );

    // Connections for Dual-Port RAM
    assign ram_data_addr = decoded_immediate_operand; // Data address is always the immediate operand
    assign ram_data_in_data = {8'h00, acc_out};      // Data to write to RAM from Accumulator


    // 3. Instruction Register (IR) / Decoder
    // The instruction_in for ir_decoder now comes from the instruction port of RAM
    // The ram_we is now ram_we_data, and ram_addr_mux_sel is no longer needed
    ir_decoder u_ir_decoder (
        .clk(clk_50mhz),
        .reset_n(key0_n),
        .instruction_in(instruction_from_ram_inst), // Instruction from RAM's Port A

        .pc_load_en(pc_load_en),
        .jump_addr(jump_addr),

        .ram_we(ram_we_data),                      // Now controls Port B's write enable
        // .ram_addr_mux_sel(ram_addr_mux_sel),    // REMOVED: No longer needed for muxing RAM address

        .alu_opcode(alu_opcode),
        .alu_a_mux_sel(alu_a_mux_sel),
        .alu_b_mux_sel(alu_b_mux_sel),

        .acc_load_en(acc_load_en),

        .immediate_operand(decoded_immediate_operand),
        .serial_out_en(serial_out_en),
        .decoded_opcode_out(decoded_opcode)
    );

    // 4. Accumulator
    accumulator u_acc (
        .clk(clk_50mhz),
        .reset_n(key0_n),
        .acc_load_en(acc_load_en),
        .data_in(acc_data_in_muxed),
        .acc_out(acc_out)
    );

    // Mux for Accumulator Data Input: Selects source for ACC loading
    // Now, data from memory operations comes from data_from_ram_data (Port B)
    assign acc_data_in_muxed =
        (decoded_opcode == OP_LOAD_ACC_IMM)  ? decoded_immediate_operand :
        (decoded_opcode == OP_LOAD_ACC_MEM)  ? data_from_ram_data[7:0]   : // Data from RAM Port B
        alu_result;

    // 5. ALU
    alu u_alu (
        .a(alu_a_input),
        .b(alu_b_input),
        .opcode(alu_opcode),
        .result(alu_result),
        .carry_out(alu_carry_out)
    );

    // Mux for ALU Operand A: In this simple CPU, ALU A is always from Accumulator
    assign alu_a_input = acc_out;

    // Mux for ALU Operand B: Selects between Immediate_Operand and Lower 8 bits of RAM data (from Port B)
    assign alu_b_input = (alu_b_mux_sel == 1'b0) ? decoded_immediate_operand : data_from_ram_data[7:0]; // Data from RAM Port B


    // --- 偵錯輸出連接 ---
    assign debug_output_acc = acc_out;
    assign debug_pc_out = pc_out;
    assign debug_instruction_out = instruction_from_ram_inst; // Now specifically instruction from Port A

endmodule